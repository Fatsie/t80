F3
3E
45
32
A0
00
00
76

